version https://git-lfs.github.com/spec/v1
oid sha256:c8cef0ee212b692a163e80bf4eda5e0a09304b9c3aa6f2b123e1553de311878b
size 104858112
